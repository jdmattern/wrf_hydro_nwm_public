netcdf \2019-08-18_00.60min.CCHC1.RFCTimeSlice {
dimensions:
	stationIdStrLen = 5 ;
	timeStrLen = 19 ;
	forecastInd = UNLIMITED ; // (289 currently)
	nseries = 1 ;
	zero = UNLIMITED ; // (0 currently)
variables:
	char stationId(stationIdStrLen) ;
		stationId:long_name = "RFC station identifer of length 5" ;
		stationId:units = "-" ;
	char issueTimeUTC(nseries, timeStrLen) ;
		issueTimeUTC:long_name = "YYYY-MM-DD_HH:mm:ss UTC" ;
		issueTimeUTC:unts = "UTC" ;
	float discharges(nseries, forecastInd) ;
		discharges:long_name = "Discharge.cubic_meters_per_second" ;
		discharges:units = "m^3/s" ;
	byte synthetic_values(nseries, forecastInd) ;
		synthetic_values:long_name = "Whether the discharge value is synthetic or orginal, 1 - synthetic, 0 - original" ;
		synthetic_values:units = "-" ;
	short totalCounts(nseries) ;
		totalCounts:long_name = "Count of forecast values" ;
		totalCounts:units = "-" ;
	short observedCounts(nseries) ;
		observedCounts:long_name = "Total observed values before T0." ;
		observedCounts:units = "-" ;
	int timeSteps(nseries) ;
		timeSteps:long_name = "Frequency/temporal resolution of forecast values" ;
		timeSteps:units = "seconds" ;
	short discharge_qualities(nseries) ;
		discharge_qualities:long_name = "Discharge quality 0 to 100 to be scaled by 100." ;
		discharge_qualities:units = "-" ;
		discharge_qualities:multfactor = "0.01" ;
	int64 queryTime(nseries) ;
		queryTime:units = "seconds since 1970-01-01 00:00:00 local TZ" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1.1|hdf5libversion=1.8.18" ;
		:fileUpdateTimeUTC = "2019-12-17_13:33:00" ;
		:sliceStartTimeUTC = "2019-12-15_00:00:00" ;
		:sliceTimeResolutionMinutes = "60" ;
		:missingValue = "-999" ;
		:newest_forecast = "0" ;
		:NWM_version_number = "v2.1" ;
data:

 stationId = "CCHC1" ;

 issueTimeUTC =
  // issueTimeUTC(0, 0-18)
    "2019-12-17_00:00:00" ;

 discharges =
  {// discharges(0, 0-288)
    0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9, 1, 1.1, 1.2, 1.3, 1.4, 1.5, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 5.1, 5.2, 5.3, 5.4, 5.5, 5.6, 5.7, 5.8, 
    5.9, 6, 6.1, 6.2, 6.3, 6.4, 6.5, 6.6, 6.7, 6.8, 6.9, 7, 7.1, 7.2, 7.3, 
    7.4, 7.5, 7.6, 7.7, 7.8, 7.9, 8, 8.1, 8.2, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 3.1, 3.2, 3.3, 3.4, 3.5, 3.6, 3.7, 3.8, 3.9, 4, 
    4.1, 4.2, 4.3, 4.4, 4.5, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 53.25485, 52.25485, 51.25485, 
    50.25485, 49.25485, 48.25485, 47.25485, 46.25485, 45.25485, 44.25485, 
    43.25485, 42.25485, 42.25485, 40.25485, 39.25485, 38.25485, 37.25485, 
    36.25485, 35.25485, 34.25485, 33.25485, 32.25485, 31.25485, 30.25485, 
    29.25485, 28.25485, 27.25485, 26.25485, 25.25485, 24.25485, 23.25485, 
    22.25485, 21.25485, 20.25485, 19.25485, 18.25485, 17.25485, 16.25485, 
    15.25485, 14.25485, 13.25485, 12.25485, 11.25485, 10.25485, 9.254851, 
    8.254851, 7.254852, 6.254852, 5.254852, 4.254852} ;

 synthetic_values =
  {// synthetic_values(0, 0-288)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0} ;

 totalCounts = 289 ;

 observedCounts = 0 ;

 timeSteps = 3600 ;

 discharge_qualities = 100 ;

 queryTime = 1576540800 ;
}
