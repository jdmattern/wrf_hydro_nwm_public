netcdf \2019-08-18_00.60min.CCHC1.RFCTimeSlice {
dimensions:
	stationIdStrLen = 5 ;
	timeStrLen = 19 ;
	forecastInd = UNLIMITED ; // (289 currently)
	nseries = 1 ;
	zero = UNLIMITED ; // (0 currently)
variables:
	char stationId(stationIdStrLen) ;
		stationId:long_name = "RFC station identifer of length 5" ;
		stationId:units = "-" ;
	char issueTimeUTC(nseries, timeStrLen) ;
		issueTimeUTC:long_name = "YYYY-MM-DD_HH:mm:ss UTC" ;
		issueTimeUTC:unts = "UTC" ;
	float discharges(nseries, forecastInd) ;
		discharges:long_name = "Discharge.cubic_meters_per_second" ;
		discharges:units = "m^3/s" ;
	byte synthetic_values(nseries, forecastInd) ;
		synthetic_values:long_name = "Whether the discharge value is synthetic or orginal, 1 - synthetic, 0 - original" ;
		synthetic_values:units = "-" ;
	short forecastCounts(nseries) ;
		forecastCounts:long_name = "Count of forecast values" ;
		forecastCounts:units = "-" ;
	int timeSteps(nseries) ;
		timeSteps:long_name = "Frequency/temporal resolution of forecast values" ;
		timeSteps:units = "seconds" ;
	short discharge_qualities(nseries) ;
		discharge_qualities:long_name = "Discharge quality 0 to 100 to be scaled by 100." ;
		discharge_qualities:units = "-" ;
		discharge_qualities:multfactor = "0.01" ;
	int64 queryTime(nseries) ;
		queryTime:units = "seconds since 1970-01-01 00:00:00 local TZ" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1.1|hdf5libversion=1.8.18" ;
		:fileUpdateTimeUTC = "2019-12-17_13:33:00" ;
		:sliceStartTimeUTC = "2019-12-15_00:00:00" ;
		:sliceTimeResolutionMinutes = "60" ;
		:missingValue = "-999" ;
		:newest_forecast = "0" ;
		:NWM_version_number = "v2.1" ;
data:

 stationId = "CCHC1" ;

 issueTimeUTC =
  // issueTimeUTC(0, 0-18)
    "2019-12-17_00:00:00" ;

 discharges =
  {// discharges(0, 0-288)
    0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9, 1, 1.1, 1.2, 1.3, 1.4, 1.5, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 5.1, 5.2, 5.3, 5.4, 5.5, 5.6, 5.7, 5.8, 
    5.9, 6, 6.1, 6.2, 6.3, 6.4, 6.5, 6.6, 6.7, 6.8, 6.9, 7.0, 
    7.1, 7.2, 7.3, 7.4, 7.5, 7.6, 
    7.7, 7.8, 7.9, 8.0, 8.1, 8.2, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 3.1, 3.2, 3.3, 3.4, 3.5, 3.6, 
    3.7, 3.8, 3.9, 4, 4.1, 4.2, 4.3, 4.4, 4.5, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 0.2548516, 
    53.2548516, 52.2548516, 51.2548516, 50.2548516, 49.2548516, 48.2548516, 
    47.2548516, 46.2548516, 45.2548516, 44.2548516, 43.2548516, 42.2548516, 
    42.2548516, 40.2548516, 39.2548516, 38.2548516, 37.2548516, 36.2548516, 
    35.2548516, 34.2548516, 33.2548516, 32.2548516, 31.2548516, 30.2548516, 
    29.2548516, 28.2548516, 27.2548516, 26.2548516, 25.2548516, 24.2548516, 
    23.2548516, 22.2548516, 21.2548516, 20.2548516, 19.2548516, 18.2548516, 
    17.2548516, 16.2548516, 15.2548516, 14.2548516, 13.2548516, 12.2548516, 
    11.2548516, 10.2548516, 9.2548516, 8.2548516, 7.2548516, 6.2548516, 
    5.2548516, 4.2548516} ;

 synthetic_values =
  {// synthetic_values(0, 0-288)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0} ;

 forecastCounts = 289 ;

 timeSteps = 3600 ;

 discharge_qualities = 100 ;

 queryTime = 1576540800 ;
}
